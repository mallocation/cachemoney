library ieee;
use ieee.std_logic_1164.all;

entity HazardDetectionUnit is
	port (
		Instruction			:	in	std_logic_vector(31 downto 0);
		RegDestFromEXStage	:	in std_logic_vector(4 downto 0);
		MEMRd_WBWr_From_EX	:	in std_logic;
		RegDestFromMEMStage	:	in 	std_logic_vector(4 downto 0);
		MEMRd_WBWr_From_MEM	:	in 	std_logic;
		RegDestFromWBStage	:	in	std_logic_vector(4 downto 0);
		WBWr_From_WB		:	in 	std_logic;
		MemReadFromEXStage  :   in std_logic;		
		HDUBranchHazards	:	out std_logic;
		HDULoadWordHazards	:	out std_logic
	);	
end HazardDetectionUnit;

architecture behavior of HazardDetectionUnit is
	signal opcode	:	std_logic_vector(2 downto 0);
	signal InstructionRD	:	std_logic_vector(4 downto 0);
	signal InstructionRS	:	std_logic_vector(4 downto 0);
	signal InstructionRT    :   std_logic_vector(4 downto 0);
begin
	opcode <= Instruction(31 downto 29);
	InstructionRD <= Instruction(28 downto 24);
	InstructionRS <= Instruction(23 downto 19);
	InstructionRT <= Instruction(18 downto 14);
	
	process(opcode, InstructionRD, InstructionRS, InstructionRT, RegDestFromEXStage, RegDestFromMEMStage, RegDestFromWBStage, MemReadFromEXStage, MEMRd_WBWr_From_EX, MEMRd_WBWr_From_MEM,WBWr_From_WB)
	begin
		HDUBranchHazards <= '0';
		HDULoadWordHazards <= '0';
		if MemReadFromEXStage = '1' and ((RegDestFromEXStage = InstructionRS) or (RegDestFromEXStage = InstructionRT)) then
			HDULoadWordHazards <= '1';
		end if;

		if opcode = "101" or opcode = "110" then -- Branch on equal, branch on not equal
			if (((InstructionRD = RegDestFromEXStage or InstructionRS = RegDestFromEXStage) and MemRD_WBWr_From_EX = '1') or
				((InstructionRD = RegDestFromMEMStage or InstructionRS = RegDestFromMEMStage) and MemRD_WBWr_From_MEM = '1') or 
				((InstructionRD = RegDestFromWBStage or InstructionRS = RegDestFromWBStage) and WBWr_From_WB = '1')) then
				HDUBranchHazards <= '1';
			else
				HDUBranchHazards <= '0';					
			end if;
		end if;
	end process;
end behavior;